module Neuronen (
input wire x 
output reg [19:0] neuronen
);
    
    reg [19:0] neuronen = 20'd0;

endmodule