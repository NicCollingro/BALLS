module sqrt(
  input  wire[14:0] in,
  output wire[9:0] out
);

  assign out =   (in >= 1024) ? 32
               : (in >= 961) ? 31
               : (in >= 900) ? 30
               : (in >= 841) ? 29
               : (in >= 784) ? 28
               : (in >= 729) ? 27
               : (in >= 676) ? 26
               : (in >= 625) ? 25
               : (in >= 576) ? 24
               : (in >= 529) ? 23
               : (in >= 484) ? 22
               : (in >= 441) ? 21
               : (in >= 400) ? 20
               : (in >= 361) ? 19
               : (in >= 324) ? 18
               : (in >= 289) ? 17
               : (in >= 256) ? 16
               : (in >= 225) ? 15
               : (in >= 196) ? 14
               : (in >= 169) ? 13
               : (in >= 144) ? 12
               : (in >= 121) ? 11
               : (in >= 100) ? 10
               : (in >=  81) ?  9
               : (in >=  64) ?  8
               : (in >=  49) ?  7
               : (in >=  36) ?  6
               : (in >=  25) ?  5
               : (in >=  16) ?  4
               : (in >=   9) ?  3
               : (in >=   4) ?  2
               : (in >=   1) ?  1
               : 0;
endmodule
